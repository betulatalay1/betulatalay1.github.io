*** SPICE deck for cell 8BitALU{sch} from library 8Bit_ALU
*** Created on Çar Ara 31, 2025 15:04:01
*** Last revised on Per Oca 01, 2026 20:55:36
*** Written on Per Oca 01, 2026 21:04:43 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SingleInverter_forFA__Inv FROM CELL SingleInverter_forFA:Inv{sch}
.SUBCKT SingleInverter_forFA__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=3U
.ENDS SingleInverter_forFA__Inv

*** SUBCIRCUIT NandGate_forFA__NAND FROM CELL NandGate_forFA:NAND{sch}
.SUBCKT NandGate_forFA__NAND A AB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AB A net@5 gnd N L=0.6U W=3U
Mnmos@1 net@5 B gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A AB vdd P L=0.6U W=3U
Mpmos@1 vdd B AB vdd P L=0.6U W=3U
.ENDS NandGate_forFA__NAND

*** SUBCIRCUIT XorGate_forFA__XOR FROM CELL XorGate_forFA:XOR{sch}
.SUBCKT XorGate_forFA__XOR A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A net@15 gnd N L=0.6U W=3U
Mnmos@1 out net@51 net@15 gnd N L=0.6U W=3U
Mnmos@2 net@15 B gnd gnd N L=0.6U W=3U
Mnmos@3 net@15 net@50 gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A net@2 vdd P L=0.6U W=3U
Mpmos@1 net@2 net@51 out vdd P L=0.6U W=3U
Mpmos@3 vdd B net@3 vdd P L=0.6U W=3U
Mpmos@4 net@3 net@50 out vdd P L=0.6U W=3U
XInv@0 A net@50 SingleInverter_forFA__Inv
XInv@1 B net@51 SingleInverter_forFA__Inv
.ENDS XorGate_forFA__XOR

*** SUBCIRCUIT HalfAdder__HalfAdder FROM CELL HalfAdder:HalfAdder{sch}
.SUBCKT HalfAdder__HalfAdder A B C S
** GLOBAL gnd
** GLOBAL vdd
XInv@0 net@10 C SingleInverter_forFA__Inv
XNAND@0 A net@10 B NandGate_forFA__NAND
XXOR@1 A B S XorGate_forFA__XOR
.ENDS HalfAdder__HalfAdder

*** SUBCIRCUIT NorGate_forFA__NOR FROM CELL NorGate_forFA:NOR{sch}
.SUBCKT NorGate_forFA__NOR A AorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AorB B gnd gnd N L=0.6U W=3U
Mnmos@1 AorB A gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A net@1 vdd P L=0.6U W=3U
Mpmos@1 net@1 B AorB vdd P L=0.6U W=3U
.ENDS NorGate_forFA__NOR

*** SUBCIRCUIT FullAdder__FullAdder FROM CELL FullAdder:FullAdder{sch}
.SUBCKT FullAdder__FullAdder A B Cin Cout S
** GLOBAL gnd
** GLOBAL vdd
XHalfAdde@0 A B net@6 net@4 HalfAdder__HalfAdder
XHalfAdde@1 Cin net@4 net@7 S HalfAdder__HalfAdder
XInv@0 net@0 Cout SingleInverter_forFA__Inv
XNOR@0 net@7 net@0 net@6 NorGate_forFA__NOR
.ENDS FullAdder__FullAdder

*** SUBCIRCUIT _8Bit_Adder__8Bit_Adder FROM CELL 8Bit_Adder:8Bit_Adder{sch}
.SUBCKT _8Bit_Adder__8Bit_Adder A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cin Cout S0 S1 S2 S3 S4 S5 S6 S7
** GLOBAL gnd
** GLOBAL vdd
XFullAdde@0 A0 B0 Cin net@0 S0 FullAdder__FullAdder
XFullAdde@1 A1 B1 net@0 net@21 S1 FullAdder__FullAdder
XFullAdde@2 A2 B2 net@21 net@28 S2 FullAdder__FullAdder
XFullAdde@3 A3 B3 net@28 net@35 S3 FullAdder__FullAdder
XFullAdde@4 A4 B4 net@35 net@42 S4 FullAdder__FullAdder
XFullAdde@5 A5 B5 net@42 net@49 S5 FullAdder__FullAdder
XFullAdde@6 A6 B6 net@49 net@56 S6 FullAdder__FullAdder
XFullAdde@7 A7 B7 net@56 Cout S7 FullAdder__FullAdder
.ENDS _8Bit_Adder__8Bit_Adder

*** SUBCIRCUIT SingleInverter_for8__Inv FROM CELL SingleInverter_for8:Inv{sch}
.SUBCKT SingleInverter_for8__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=3U
.ENDS SingleInverter_for8__Inv

*** SUBCIRCUIT _8Bit_Inv__8Bit_Inv FROM CELL 8Bit_Inv:8Bit_Inv{sch}
.SUBCKT _8Bit_Inv__8Bit_Inv A0 A0not A1 A1not A2 A2not A3 A3not A4 A4not A5 A5not A6 A6not A7 A7not
** GLOBAL gnd
** GLOBAL vdd
XInv@0 A0 A0not SingleInverter_for8__Inv
XInv@1 A1 A1not SingleInverter_for8__Inv
XInv@2 A2 A2not SingleInverter_for8__Inv
XInv@3 A3 A3not SingleInverter_for8__Inv
XInv@4 A4 A4not SingleInverter_for8__Inv
XInv@5 A5 A5not SingleInverter_for8__Inv
XInv@6 A6 A6not SingleInverter_for8__Inv
XInv@7 A7 A7not SingleInverter_for8__Inv
.ENDS _8Bit_Inv__8Bit_Inv

*** SUBCIRCUIT _8Bit_SUB__8Bit_SUB FROM CELL 8Bit_SUB:8Bit_SUB{sch}
.SUBCKT _8Bit_SUB__8Bit_SUB A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cout Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
X_8Bit_Add@0 A0 A1 A2 A3 A4 A5 A6 A7 net@9 net@11 net@14 net@17 net@20 net@23 net@26 net@29 vdd Cout Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 _8Bit_Adder__8Bit_Adder
X_8Bit_Inv@0 B0 net@9 B1 net@11 B2 net@14 B3 net@17 B4 net@20 B5 net@23 B6 net@26 B7 net@29 _8Bit_Inv__8Bit_Inv
.ENDS _8Bit_SUB__8Bit_SUB

*** SUBCIRCUIT Inverter_forZERO__Inv FROM CELL Inverter_forZERO:Inv{sch}
.SUBCKT Inverter_forZERO__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=3U
.ENDS Inverter_forZERO__Inv

*** SUBCIRCUIT NorGate_forZERO__NOR FROM CELL NorGate_forZERO:NOR{sch}
.SUBCKT NorGate_forZERO__NOR A AorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AorB B gnd gnd N L=0.6U W=3U
Mnmos@1 AorB A gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A net@1 vdd P L=0.6U W=3U
Mpmos@1 net@1 B AorB vdd P L=0.6U W=3U
.ENDS NorGate_forZERO__NOR

*** SUBCIRCUIT OrGate__or FROM CELL OrGate:or{sch}
.SUBCKT OrGate__or A B out
** GLOBAL gnd
** GLOBAL vdd
XInv@0 net@0 out Inverter_forZERO__Inv
XNOR@0 A net@0 B NorGate_forZERO__NOR
.ENDS OrGate__or

*** SUBCIRCUIT zeroflag__zeroflag FROM CELL zeroflag:zeroflag{sch}
.SUBCKT zeroflag__zeroflag A0 A1 A2 A3 A4 A5 A6 A7 out
** GLOBAL gnd
** GLOBAL vdd
XInv@7 net@192 out Inverter_forZERO__Inv
Xor@0 A0 A1 net@175 OrGate__or
Xor@1 A2 A3 net@177 OrGate__or
Xor@2 A4 A5 net@179 OrGate__or
Xor@3 A6 A7 net@181 OrGate__or
Xor@4 net@175 net@177 net@185 OrGate__or
Xor@5 net@179 net@181 net@183 OrGate__or
Xor@6 net@185 net@183 net@192 OrGate__or
.ENDS zeroflag__zeroflag

*** SUBCIRCUIT _8BitSUB_COMP__8BitSUB_COMP FROM CELL 8BitSUB_COMP:8BitSUB_COMP{sch}
.SUBCKT _8BitSUB_COMP__8BitSUB_COMP A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Equal Greater Less Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
X_8Bit_SUB@0 A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 net@16 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 _8Bit_SUB__8Bit_SUB
XInv@1 net@16 Less Inverter_forZERO__Inv
XNOR@0 Equal Greater Less NorGate_forZERO__NOR
Xzeroflag@0 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 Equal zeroflag__zeroflag
.ENDS _8BitSUB_COMP__8BitSUB_COMP

*** SUBCIRCUIT NandGate_for8NAND__NAND FROM CELL NandGate_for8NAND:NAND{sch}
.SUBCKT NandGate_for8NAND__NAND A AB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AB A net@5 gnd N L=0.6U W=3U
Mnmos@1 net@5 B gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A AB vdd P L=0.6U W=3U
Mpmos@1 vdd B AB vdd P L=0.6U W=3U
.ENDS NandGate_for8NAND__NAND

*** SUBCIRCUIT _8Bit_NAND__8Bit_NAND FROM CELL 8Bit_NAND:8Bit_NAND{sch}
.SUBCKT _8Bit_NAND__8Bit_NAND A0 A1 A2 A3 A4 A5 A6 A7 AB0 AB1 AB2 AB3 AB4 AB5 AB6 AB7 B0 B1 B2 B3 B4 B5 B6 B7
** GLOBAL gnd
** GLOBAL vdd
XNAND@0 A0 AB0 B0 NandGate_for8NAND__NAND
XNAND@1 A1 AB1 B1 NandGate_for8NAND__NAND
XNAND@2 A2 AB2 B2 NandGate_for8NAND__NAND
XNAND@3 A3 AB3 B3 NandGate_for8NAND__NAND
XNAND@4 A4 AB4 B4 NandGate_for8NAND__NAND
XNAND@5 A5 AB5 B5 NandGate_for8NAND__NAND
XNAND@6 A6 AB6 B6 NandGate_for8NAND__NAND
XNAND@7 A7 AB7 B7 NandGate_for8NAND__NAND
.ENDS _8Bit_NAND__8Bit_NAND

*** SUBCIRCUIT _8Bit_AND__8Bit_AND FROM CELL 8Bit_AND:8Bit_AND{sch}
.SUBCKT _8Bit_AND__8Bit_AND A0 A1 A2 A3 A4 A5 A6 A7 AandB0 AandB1 AandB2 AandB3 AandB4 AandB5 AandB6 AandB7 B0 B1 B2 B3 B4 B5 B6 B7
** GLOBAL gnd
** GLOBAL vdd
X_8Bit_Inv@0 net@0 AandB0 net@2 AandB1 net@5 AandB2 net@13 AandB3 net@16 AandB4 net@19 AandB5 net@24 AandB6 net@22 AandB7 _8Bit_Inv__8Bit_Inv
X_8Bit_NAN@0 A0 A1 A2 A3 A4 A5 A6 A7 net@0 net@2 net@5 net@13 net@16 net@19 net@24 net@22 B0 B1 B2 B3 B4 B5 B6 B7 _8Bit_NAND__8Bit_NAND
.ENDS _8Bit_AND__8Bit_AND

*** SUBCIRCUIT NorGate_for8NOR__NOR FROM CELL NorGate_for8NOR:NOR{sch}
.SUBCKT NorGate_for8NOR__NOR A AorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AorB B gnd gnd N L=0.6U W=3U
Mnmos@1 AorB A gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A net@1 vdd P L=0.6U W=3U
Mpmos@1 net@1 B AorB vdd P L=0.6U W=3U
.ENDS NorGate_for8NOR__NOR

*** SUBCIRCUIT _8Bit_NOR__8Bit_NOR FROM CELL 8Bit_NOR:8Bit_NOR{sch}
.SUBCKT _8Bit_NOR__8Bit_NOR A0 A1 A2 A3 A4 A5 A6 A7 AorB0 AorB1 AorB2 AorB3 AorB4 AorB5 AorB6 AorB7 B0 B1 B2 B3 B4 B5 B6 B7
** GLOBAL gnd
** GLOBAL vdd
XNOR@0 A0 AorB0 B0 NorGate_for8NOR__NOR
XNOR@1 A1 AorB1 B1 NorGate_for8NOR__NOR
XNOR@2 A2 AorB2 B2 NorGate_for8NOR__NOR
XNOR@3 A3 AorB3 B3 NorGate_for8NOR__NOR
XNOR@4 A4 AorB4 B4 NorGate_for8NOR__NOR
XNOR@5 A5 AorB5 B5 NorGate_for8NOR__NOR
XNOR@6 A6 AorB6 B6 NorGate_for8NOR__NOR
XNOR@7 A7 AorB7 B7 NorGate_for8NOR__NOR
.ENDS _8Bit_NOR__8Bit_NOR

*** SUBCIRCUIT _8Bit_OR__8Bit_OR FROM CELL 8Bit_OR:8Bit_OR{sch}
.SUBCKT _8Bit_OR__8Bit_OR A0 A1 A2 A3 A4 A5 A6 A7 AorB0 AorB1 AorB2 AorB3 AorB4 AorB5 AorB6 AorB7 B0 B1 B2 B3 B4 B5 B6 B7
** GLOBAL gnd
** GLOBAL vdd
X_8Bit_Inv@0 net@0 AorB0 net@2 AorB1 net@4 AorB2 net@6 AorB3 net@8 AorB4 net@10 AorB5 net@13 AorB6 net@16 AorB7 _8Bit_Inv__8Bit_Inv
X_8Bit_NOR@0 A0 A1 A2 A3 A4 A5 A6 A7 net@0 net@2 net@4 net@6 net@8 net@10 net@13 net@16 B0 B1 B2 B3 B4 B5 B6 B7 _8Bit_NOR__8Bit_NOR
.ENDS _8Bit_OR__8Bit_OR

*** SUBCIRCUIT SingleInverter_for8XOR__Inv FROM CELL SingleInverter_for8XOR:Inv{sch}
.SUBCKT SingleInverter_for8XOR__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=3U
.ENDS SingleInverter_for8XOR__Inv

*** SUBCIRCUIT XorGate_for8XOR__XOR FROM CELL XorGate_for8XOR:XOR{sch}
.SUBCKT XorGate_for8XOR__XOR A B out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out A net@15 gnd N L=0.6U W=3U
Mnmos@1 out net@51 net@15 gnd N L=0.6U W=3U
Mnmos@2 net@15 B gnd gnd N L=0.6U W=3U
Mnmos@3 net@15 net@50 gnd gnd N L=0.6U W=3U
Mpmos@0 vdd A net@2 vdd P L=0.6U W=3U
Mpmos@1 net@2 net@51 out vdd P L=0.6U W=3U
Mpmos@3 vdd B net@3 vdd P L=0.6U W=3U
Mpmos@4 net@3 net@50 out vdd P L=0.6U W=3U
XInv@0 A net@50 SingleInverter_for8XOR__Inv
XInv@1 B net@51 SingleInverter_for8XOR__Inv
.ENDS XorGate_for8XOR__XOR

*** SUBCIRCUIT _8Bit_XOR__8Bit_XOR FROM CELL 8Bit_XOR:8Bit_XOR{sch}
.SUBCKT _8Bit_XOR__8Bit_XOR A0 A1 A2 A3 A4 A5 A6 A7 AxorB_0 AxorB_1 AxorB_2 AxorB_3 AxorB_4 AxorB_5 AxorB_6 AxorB_7 B0 B1 B2 B3 B4 B5 B6 B7
** GLOBAL gnd
** GLOBAL vdd
XXOR@0 A0 B0 AxorB_0 XorGate_for8XOR__XOR
XXOR@1 A1 B1 AxorB_1 XorGate_for8XOR__XOR
XXOR@2 A2 B2 AxorB_2 XorGate_for8XOR__XOR
XXOR@3 A3 B3 AxorB_3 XorGate_for8XOR__XOR
XXOR@4 A4 B4 AxorB_4 XorGate_for8XOR__XOR
XXOR@5 A5 B5 AxorB_5 XorGate_for8XOR__XOR
XXOR@6 A6 B6 AxorB_6 XorGate_for8XOR__XOR
XXOR@7 A7 B7 AxorB_7 XorGate_for8XOR__XOR
.ENDS _8Bit_XOR__8Bit_XOR

*** SUBCIRCUIT SingleInverter_for16MUX__Inv FROM CELL SingleInverter_for16MUX:Inv{sch}
.SUBCKT SingleInverter_for16MUX__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=3U
.ENDS SingleInverter_for16MUX__Inv

*** SUBCIRCUIT MUX2_1__MUX2_1 FROM CELL MUX2_1:MUX2_1{sch}
.SUBCKT MUX2_1__MUX2_1 A B out S
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 A net@22 out gnd N L=0.6U W=3U
Mnmos@1 B S out gnd N L=0.6U W=3U
Mpmos@0 out S A vdd P L=0.6U W=3U
Mpmos@1 out net@22 B vdd P L=0.6U W=3U
XInv@1 S net@22 SingleInverter_for16MUX__Inv
.ENDS MUX2_1__MUX2_1

*** SUBCIRCUIT MUX4_1__MUX4_1 FROM CELL MUX4_1:MUX4_1{sch}
.SUBCKT MUX4_1__MUX4_1 out S0 S1 I0 I1 I2 I3
** GLOBAL gnd
** GLOBAL vdd
XMUX2_1@0 I2 I3 net@16 S0 MUX2_1__MUX2_1
XMUX2_1@1 I0 I1 net@13 S0 MUX2_1__MUX2_1
XMUX2_1@2 net@13 net@16 out S1 MUX2_1__MUX2_1
.ENDS MUX4_1__MUX4_1

*** SUBCIRCUIT MUX16_1__MUX16_1 FROM CELL MUX16_1:MUX16_1{sch}
.SUBCKT MUX16_1__MUX16_1 out S0 S1 S2 S3 I0 I1 I10 I11 I12 I13 I14 I15 I2 I3 I4 I5 I6 I7 I8 I9
** GLOBAL gnd
** GLOBAL vdd
XMUX4_1@0 net@0 S0 S1 I0 I1 I2 I3 MUX4_1__MUX4_1
XMUX4_1@1 net@3 S0 S1 I4 I5 I6 I7 MUX4_1__MUX4_1
XMUX4_1@2 net@6 S0 S1 I8 I9 I10 I11 MUX4_1__MUX4_1
XMUX4_1@3 net@13 S0 S1 I12 I13 I14 I15 MUX4_1__MUX4_1
XMUX4_1@4 out S2 S3 net@0 net@3 net@6 net@13 MUX4_1__MUX4_1
.ENDS MUX16_1__MUX16_1

*** SUBCIRCUIT Inverter_aleft__Inv FROM CELL Inverter_aleft:Inv{sch}
.SUBCKT Inverter_aleft__Inv in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd N L=0.6U W=3U
Mpmos@0 vdd in out vdd P L=0.6U W=3U
.ENDS Inverter_aleft__Inv

*** SUBCIRCUIT _8Bit_Inv_aleft__8Bit_Inv FROM CELL 8Bit_Inv_aleft:8Bit_Inv{sch}
.SUBCKT _8Bit_Inv_aleft__8Bit_Inv A0 A1 A2 A3 A4 A5 A6 A7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
XInv@0 A0 Y0 Inverter_aleft__Inv
XInv@1 A1 Y1 Inverter_aleft__Inv
XInv@2 A2 Y2 Inverter_aleft__Inv
XInv@3 A3 Y3 Inverter_aleft__Inv
XInv@4 A4 Y4 Inverter_aleft__Inv
XInv@5 A5 Y5 Inverter_aleft__Inv
XInv@6 A6 Y6 Inverter_aleft__Inv
XInv@7 A7 Y7 Inverter_aleft__Inv
.ENDS _8Bit_Inv_aleft__8Bit_Inv

*** SUBCIRCUIT buf_8__buf_8 FROM CELL buf_8:buf_8{sch}
.SUBCKT buf_8__buf_8 A0 A1 A2 A3 A4 A5 A6 A7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
X_8Bit_Inv@0 A0 A1 A2 A3 A4 A5 A6 A7 net@0 net@1 net@2 net@3 net@4 net@5 net@6 net@7 _8Bit_Inv_aleft__8Bit_Inv
X_8Bit_Inv@1 net@0 net@1 net@2 net@3 net@4 net@5 net@6 net@7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 _8Bit_Inv_aleft__8Bit_Inv
.ENDS buf_8__buf_8

*** SUBCIRCUIT a_left_shift__a_left_shift FROM CELL a_left_shift:a_left_shift{sch}
.SUBCKT a_left_shift__a_left_shift in0 in1 in2 in3 in4 in5 in6 in7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
Xbuf_8@0 gnd in0 in1 in2 in3 in4 in5 in6 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 buf_8__buf_8
.ENDS a_left_shift__a_left_shift

*** SUBCIRCUIT a_right_shift__a_right_shift FROM CELL a_right_shift:a_right_shift{sch}
.SUBCKT a_right_shift__a_right_shift in0 in1 in2 in3 in4 in5 in6 in7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
Xbuf_8@0 in1 in2 in3 in4 in5 in6 gnd in7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 buf_8__buf_8
.ENDS a_right_shift__a_right_shift

*** SUBCIRCUIT left_shift__left_shift FROM CELL left_shift:left_shift{sch}
.SUBCKT left_shift__left_shift in0 in1 in2 in3 in4 in5 in6 in7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
Xbuf_8@0 gnd in0 in1 in2 in3 in4 in5 in6 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 buf_8__buf_8
.ENDS left_shift__left_shift

*** SUBCIRCUIT right_shift__right_shift FROM CELL right_shift:right_shift{sch}
.SUBCKT right_shift__right_shift in0 in1 in2 in3 in4 in5 in6 in7 Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
** GLOBAL gnd
** GLOBAL vdd
Xbuf_8@0 in1 in2 in3 in4 in5 in6 in7 gnd Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 buf_8__buf_8
.ENDS right_shift__right_shift

.global gnd vdd

*** TOP LEVEL CELL: 8BitALU{sch}
X_8BitSUB_@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 net@182 net@185 net@188 net@177 net@150 net@153 net@158 net@163 net@166 net@169 net@172 _8BitSUB_COMP__8BitSUB_COMP
X_8Bit_AND@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@191 net@194 net@198 net@201 net@207 net@212 net@215 net@220 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 _8Bit_AND__8Bit_AND
X_8Bit_Add@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 gnd Cout net@113 net@117 net@120 net@124 net@128 net@132 net@137 net@140 _8Bit_Adder__8Bit_Adder
X_8Bit_Inv@0 net@624 net@297 net@625 net@302 net@628 net@305 net@631 net@310 net@633 net@315 net@730 net@320 net@637 net@325 net@796 net@328 _8Bit_Inv__8Bit_Inv
X_8Bit_NAN@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@409 net@428 net@433 net@438 net@444 net@449 net@454 net@457 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 _8Bit_NAND__8Bit_NAND
X_8Bit_NOR@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@465 net@472 net@478 net@483 net@488 net@493 net@498 net@510 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 _8Bit_NOR__8Bit_NOR
X_8Bit_OR@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@225 net@228 net@231 net@236 net@239 net@244 net@249 net@254 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 _8Bit_OR__8Bit_OR
X_8Bit_XOR@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@259 net@264 net@267 net@275 net@279 net@282 net@287 net@292 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 _8Bit_XOR__8Bit_XOR
XMUX16_1@0 Result0 S0 S1 S2 S3 net@113 net@177 net@185 net@188 net@409 net@465 net@514 net@569 net@191 net@225 net@259 net@297 net@334 net@372 MUX16_1@0_I8 net@182 MUX16_1__MUX16_1
XMUX16_1@1 Result1 S0 S1 S2 S3 net@117 net@150 gnd gnd net@428 net@472 net@521 net@577 net@194 net@228 net@264 net@302 net@339 net@377 MUX16_1@1_I8 gnd MUX16_1__MUX16_1
XMUX16_1@2 Result2 S0 S1 S2 S3 net@120 net@153 gnd gnd net@433 net@478 net@526 net@584 net@198 net@231 net@267 net@305 net@344 net@382 MUX16_1@2_I8 gnd MUX16_1__MUX16_1
XMUX16_1@3 Result3 S0 S1 S2 S3 net@124 net@158 gnd gnd net@438 net@483 net@531 net@589 net@201 net@236 net@275 net@310 net@349 net@387 MUX16_1@3_I8 gnd MUX16_1__MUX16_1
XMUX16_1@4 Result4 S0 S1 S2 S3 net@128 net@163 gnd gnd net@444 net@488 net@536 net@602 net@207 net@239 net@279 net@315 net@358 net@393 MUX16_1@4_I8 gnd MUX16_1__MUX16_1
XMUX16_1@5 Result5 S0 S1 S2 S3 net@132 net@166 gnd gnd net@449 net@493 net@543 net@607 net@212 net@244 net@282 net@320 net@361 net@397 MUX16_1@5_I8 gnd MUX16_1__MUX16_1
XMUX16_1@6 Result6 S0 S1 S2 S3 net@137 net@169 gnd gnd net@454 net@498 net@553 net@612 net@215 net@249 net@287 net@325 net@366 net@401 MUX16_1@6_I8 gnd MUX16_1__MUX16_1
XMUX16_1@7 Result7 S0 S1 S2 S3 net@140 net@172 gnd gnd net@457 net@510 net@564 net@617 net@220 net@254 net@292 net@328 net@369 net@406 MUX16_1@7_I8 gnd MUX16_1__MUX16_1
Xa_left_s@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@514 net@521 net@526 net@531 net@536 net@543 net@553 net@564 a_left_shift__a_left_shift
Xa_right_@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@569 net@577 net@584 net@589 net@602 net@607 net@612 net@617 a_right_shift__a_right_shift
Xbuf_8@0 A0 A1 A2 A3 A4 A5 A6 A7 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 buf_8__buf_8
Xbuf_8@1 B0 B1 B2 B3 B4 B5 B6 B7 net@1039 net@1042 net@1045 net@1050 net@1053 net@1056 net@1059 net@1062 buf_8__buf_8
Xleft_shi@2 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@334 net@339 net@344 net@349 net@358 net@361 net@366 net@369 left_shift__left_shift
Xright_sh@0 net@624 net@625 net@628 net@631 net@633 net@730 net@637 net@796 net@372 net@377 net@382 net@387 net@393 net@397 net@401 net@406 right_shift__right_shift

* Spice Code nodes in cell cell '8BitALU{sch}'
vdd vdd 0 DC 5 
vS0 s0 0 DC 0
vS1 s1 0 DC 5 
vS2 s2 0 DC 5 
vS3 s3 0 DC 5 
va0 A0 0 DC pwl 10n 0 20n 0 50n 0 60n 0  
vb0 B0 0 DC pwl 10n 0 20n 5 50n 5 60n 0  
va1 A1 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb1 B1 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va2 A2 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb2 B2 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
va3 A3 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb3 B3 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va4 A4 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
vb4 B4 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va5 A5 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
vb5 B5 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va6 A6 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb6 B6 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va7 A7 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
vb7 B7 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
.tran 200n 
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
* Trailer cards described in this file:
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
.END
