*** SPICE deck for cell 8Bit_NAND{lay} from library 8Bit_NAND
*** Created on Pzt Ara 22, 2025 21:42:56
*** Last revised on Pzt Ara 22, 2025 22:11:45
*** Written on Sal Ara 23, 2025 21:28:16 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT NandGate_for8NAND__NAND FROM CELL NandGate_for8NAND:NAND{lay}
.SUBCKT NandGate_for8NAND__NAND A AB B gnd vdd
Mnmos@1 AB A net@6 gnd N L=0.6U W=3U AS=2.7P AD=5.25P PS=4.8U PD=7.5U
Mnmos@2 net@6 B gnd gnd N L=0.6U W=3U AS=20.25P AD=2.7P PS=31.5U PD=4.8U
Mpmos@0 vdd A AB vdd P L=0.6U W=3U AS=5.25P AD=13.5P PS=7.5U PD=21U
Mpmos@1 AB B vdd vdd P L=0.6U W=3U AS=13.5P AD=5.25P PS=21U PD=7.5U
.ENDS NandGate_for8NAND__NAND

*** TOP LEVEL CELL: 8Bit_NAND{lay}
XNAND@0 A0 AB0 B0 gnd vdd NandGate_for8NAND__NAND
XNAND@1 A1 AB1 B1 gnd vdd NandGate_for8NAND__NAND
XNAND@2 A2 AB2 B2 gnd vdd NandGate_for8NAND__NAND
XNAND@3 A3 AB3 B3 gnd vdd NandGate_for8NAND__NAND
XNAND@4 A4 AB4 B4 gnd vdd NandGate_for8NAND__NAND
XNAND@5 A5 AB5 B5 gnd vdd NandGate_for8NAND__NAND
XNAND@6 A6 AB6 B6 gnd vdd NandGate_for8NAND__NAND
XNAND@7 A7 AB7 B7 gnd vdd NandGate_for8NAND__NAND

* Spice Code nodes in cell cell '8Bit_NAND{lay}'
vdd vdd 0 DC 5
va0 A0 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb0 B0 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va1 A1 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb1 B1 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va2 A2 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb2 B2 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va3 A3 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb3 B3 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va4 A4 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb4 B4 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va5 A5 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb5 B5 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va6 A6 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb6 B6 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va7 A7 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb7 B7 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.tran 200n
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
* Trailer cards described in this file:
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
.END
