*** SPICE deck for cell 8Bit_SUB{lay} from library 8Bit_SUB
*** Created on Cmt Ara 27, 2025 21:41:37
*** Last revised on Cmt Ara 27, 2025 22:24:56
*** Written on Cmt Ara 27, 2025 22:24:59 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SingleInverter_forFA__Inv FROM CELL SingleInverter_forFA:Inv{lay}
.SUBCKT SingleInverter_forFA__Inv gnd in out vdd
Mnmos@0 gnd in out gnd N L=0.6U W=3U AS=6.75P AD=18P PS=10.5U PD=28.5U
Mpmos@0 vdd in out vdd P L=0.6U W=3U AS=6.75P AD=20.25P PS=10.5U PD=29.1U
.ENDS SingleInverter_forFA__Inv

*** SUBCIRCUIT NandGate_forFA__NAND FROM CELL NandGate_forFA:NAND{lay}
.SUBCKT NandGate_forFA__NAND A AB B gnd vdd
Mnmos@1 AB A net@6 gnd N L=0.6U W=3U AS=2.7P AD=5.25P PS=4.8U PD=7.5U
Mnmos@2 net@6 B gnd gnd N L=0.6U W=3U AS=20.25P AD=2.7P PS=31.5U PD=4.8U
Mpmos@0 vdd A AB vdd P L=0.6U W=3U AS=5.25P AD=13.5P PS=7.5U PD=21U
Mpmos@1 AB B vdd vdd P L=0.6U W=3U AS=13.5P AD=5.25P PS=21U PD=7.5U
.ENDS NandGate_forFA__NAND

*** SUBCIRCUIT XorGate_forFA__XOR FROM CELL XorGate_forFA:XOR{lay}
.SUBCKT XorGate_forFA__XOR A B gnd out vdd
Mnmos@0 net@6 A out gnd N L=0.6U W=3U AS=4.275P AD=5.4P PS=5.85U PD=8.1U
Mnmos@1 out net@17 net@6 gnd N L=0.6U W=3U AS=5.4P AD=4.275P PS=8.1U PD=5.85U
Mnmos@2 net@6 net@28 gnd gnd N L=0.6U W=3U AS=17.775P AD=5.4P PS=25.35U PD=8.1U
Mnmos@3 gnd B net@6 gnd N L=0.6U W=3U AS=5.4P AD=17.775P PS=8.1U PD=25.35U
Mnmos@4 gnd A net@28 gnd N L=0.6U W=3U AS=6.75P AD=17.775P PS=10.5U PD=25.35U
Mnmos@5 net@17 B gnd gnd N L=0.6U W=3U AS=17.775P AD=6.75P PS=25.35U PD=10.5U
Mpmos@0 vdd A net@1 vdd P L=0.6U W=3U AS=2.25P AD=21.6P PS=4.5U PD=27.9U
Mpmos@2 net@1 net@17 out vdd P L=0.6U W=3U AS=4.275P AD=2.25P PS=5.85U PD=4.5U
Mpmos@3 out net@28 net@4 vdd P L=0.6U W=3U AS=2.7P AD=4.275P PS=4.8U PD=5.85U
Mpmos@4 net@4 B vdd vdd P L=0.6U W=3U AS=21.6P AD=2.7P PS=27.9U PD=4.8U
Mpmos@5 vdd A net@28 vdd P L=0.6U W=3U AS=6.75P AD=21.6P PS=10.5U PD=27.9U
Mpmos@6 net@17 B vdd vdd P L=0.6U W=3U AS=21.6P AD=6.75P PS=27.9U PD=10.5U
.ENDS XorGate_forFA__XOR

*** SUBCIRCUIT HalfAdder__HalfAdder FROM CELL HalfAdder:HalfAdder{lay}
.SUBCKT HalfAdder__HalfAdder A B C gnd S vdd
XInv@0 gnd net@55 C vdd SingleInverter_forFA__Inv
XNAND@0 A net@55 B gnd vdd NandGate_forFA__NAND
XXOR@0 A B gnd S vdd XorGate_forFA__XOR
.ENDS HalfAdder__HalfAdder

*** SUBCIRCUIT NorGate_forFA__NOR FROM CELL NorGate_forFA:NOR{lay}
.SUBCKT NorGate_forFA__NOR A AorB B gnd vdd
Mnmos@0 gnd A AorB gnd N L=0.6U W=3U AS=5.25P AD=13.5P PS=7.5U PD=21U
Mnmos@1 AorB B gnd gnd N L=0.6U W=3U AS=13.5P AD=5.25P PS=21U PD=7.5U
Mpmos@0 vdd A net@6 vdd P L=0.6U W=3U AS=2.25P AD=22.95P PS=4.5U PD=32.1U
Mpmos@1 net@6 B AorB vdd P L=0.6U W=3U AS=5.25P AD=2.25P PS=7.5U PD=4.5U
.ENDS NorGate_forFA__NOR

*** SUBCIRCUIT FullAdder__FullAdder FROM CELL FullAdder:FullAdder{lay}
.SUBCKT FullAdder__FullAdder A B Cin Cout gnd S vdd
XHalfAdde@0 A B net@41 gnd net@8 vdd HalfAdder__HalfAdder
XHalfAdde@1 Cin net@8 net@46 gnd S vdd HalfAdder__HalfAdder
XInv@0 gnd net@47 Cout vdd SingleInverter_forFA__Inv
XNOR@1 net@41 net@47 net@46 gnd vdd NorGate_forFA__NOR
.ENDS FullAdder__FullAdder

*** SUBCIRCUIT _8Bit_Adder__8Bit_Adder FROM CELL 8Bit_Adder:8Bit_Adder{lay}
.SUBCKT _8Bit_Adder__8Bit_Adder A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 Cin Cout gnd S0 S1 S2 S3 S4 S5 S6 S7 vdd
XFullAdde@0 A0 B0 Cin net@80 gnd S0 vdd FullAdder__FullAdder
XFullAdde@1 A1 B1 net@80 net@88 gnd S1 vdd FullAdder__FullAdder
XFullAdde@2 A2 B2 net@88 net@99 gnd S2 vdd FullAdder__FullAdder
XFullAdde@3 A3 B3 net@99 net@110 gnd S3 vdd FullAdder__FullAdder
XFullAdde@4 A4 B4 net@110 net@118 gnd S4 vdd FullAdder__FullAdder
XFullAdde@5 A5 B5 net@118 net@124 gnd S5 vdd FullAdder__FullAdder
XFullAdde@6 A6 B6 net@124 net@134 gnd S6 vdd FullAdder__FullAdder
XFullAdde@7 A7 B7 net@134 Cout gnd S7 vdd FullAdder__FullAdder
.ENDS _8Bit_Adder__8Bit_Adder

*** SUBCIRCUIT SingleInverter_for8__Inv FROM CELL SingleInverter_for8:Inv{lay}
.SUBCKT SingleInverter_for8__Inv gnd in out vdd
Mnmos@0 gnd in out gnd N L=0.6U W=3U AS=6.75P AD=18P PS=10.5U PD=28.5U
Mpmos@0 vdd in out vdd P L=0.6U W=3U AS=6.75P AD=20.25P PS=10.5U PD=29.1U
.ENDS SingleInverter_for8__Inv

*** SUBCIRCUIT _8Bit_Inv__8Bit_Inv FROM CELL 8Bit_Inv:8Bit_Inv{lay}
.SUBCKT _8Bit_Inv__8Bit_Inv A0 A0not A1 A1not A2 A2not A3 A3not A4 A4not A5 A5not A6 A6not A7 A7not gnd vdd
XInv@0 gnd A0 A0not vdd SingleInverter_for8__Inv
XInv@1 gnd A1 A1not vdd SingleInverter_for8__Inv
XInv@2 gnd A2 A2not vdd SingleInverter_for8__Inv
XInv@3 gnd A3 A3not vdd SingleInverter_for8__Inv
XInv@4 gnd A4 A4not vdd SingleInverter_for8__Inv
XInv@5 gnd A5 A5not vdd SingleInverter_for8__Inv
XInv@6 gnd A6 A6not vdd SingleInverter_for8__Inv
XInv@7 gnd A7 A7not vdd SingleInverter_for8__Inv
.ENDS _8Bit_Inv__8Bit_Inv

*** TOP LEVEL CELL: 8Bit_SUB{lay}
X_8Bit_Add@0 A0 A1 A2 A3 A4 A5 A6 A7 net@0 net@4 net@10 net@17 net@21 net@25 net@29 net@36 vdd Cout gnd Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 vdd _8Bit_Adder__8Bit_Adder
X_8Bit_Inv@0 B0 net@0 B1 net@4 B2 net@10 B3 net@17 B4 net@21 B5 net@25 B6 net@29 B7 net@36 gnd vdd _8Bit_Inv__8Bit_Inv

* Spice Code nodes in cell cell '8Bit_SUB{lay}'
vdd vdd 0 DC 5 
va0 A0 0 DC pwl 10n 0 20n 5 50n 5 60n 0  
vb0 B0 0 DC pwl 10n 0 20n 5 50n 5 60n 0  
va1 A1 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb1 B1 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va2 A2 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
vb2 B2 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
va3 A3 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
vb3 B3 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
va4 A4 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb4 B4 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
va5 A5 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb5 B5 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va6 A6 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
vb6 B6 0 DC pwl 10n 0 20n 0 50n 0 60n 0 
va7 A7 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
vb7 B7 0 DC pwl 10n 0 20n 5 50n 5 60n 0 
.tran 200n 
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
* Trailer cards described in this file:
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
.END
