*** SPICE deck for cell 8Bit_AND{lay} from library 8Bit_AND
*** Created on Çar Ara 24, 2025 17:01:13
*** Last revised on Çar Ara 24, 2025 17:22:12
*** Written on Çar Ara 24, 2025 17:22:14 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT SingleInverter_for8__Inv FROM CELL SingleInverter_for8:Inv{lay}
.SUBCKT SingleInverter_for8__Inv gnd in out vdd
Mnmos@0 gnd in out gnd N L=0.6U W=3U AS=6.75P AD=18P PS=10.5U PD=28.5U
Mpmos@0 vdd in out vdd P L=0.6U W=3U AS=6.75P AD=20.25P PS=10.5U PD=29.1U
.ENDS SingleInverter_for8__Inv

*** SUBCIRCUIT _8Bit_Inv__8Bit_Inv FROM CELL 8Bit_Inv{lay}
.SUBCKT _8Bit_Inv__8Bit_Inv A0 A0not A1 A1not A2 A2not A3 A3not A4 A4not A5 A5not A6 A6not A7 A7not gnd vdd
XInv@0 gnd A0 A0not vdd SingleInverter_for8__Inv
XInv@1 gnd A1 A1not vdd SingleInverter_for8__Inv
XInv@2 gnd A2 A2not vdd SingleInverter_for8__Inv
XInv@3 gnd A3 A3not vdd SingleInverter_for8__Inv
XInv@4 gnd A4 A4not vdd SingleInverter_for8__Inv
XInv@5 gnd A5 A5not vdd SingleInverter_for8__Inv
XInv@6 gnd A6 A6not vdd SingleInverter_for8__Inv
XInv@7 gnd A7 A7not vdd SingleInverter_for8__Inv
.ENDS _8Bit_Inv__8Bit_Inv

*** SUBCIRCUIT NandGate_for8NAND__NAND FROM CELL NandGate_for8NAND:NAND{lay}
.SUBCKT NandGate_for8NAND__NAND A AB B gnd vdd
Mnmos@1 AB A net@6 gnd N L=0.6U W=3U AS=2.7P AD=5.25P PS=4.8U PD=7.5U
Mnmos@2 net@6 B gnd gnd N L=0.6U W=3U AS=20.25P AD=2.7P PS=31.5U PD=4.8U
Mpmos@0 vdd A AB vdd P L=0.6U W=3U AS=5.25P AD=13.5P PS=7.5U PD=21U
Mpmos@1 AB B vdd vdd P L=0.6U W=3U AS=13.5P AD=5.25P PS=21U PD=7.5U
.ENDS NandGate_for8NAND__NAND

*** SUBCIRCUIT _8Bit_NAND__8Bit_NAND FROM CELL 8Bit_NAND:8Bit_NAND{lay}
.SUBCKT _8Bit_NAND__8Bit_NAND A0 A1 A2 A3 A4 A5 A6 A7 AB0 AB1 AB2 AB3 AB4 AB5 AB6 AB7 B0 B1 B2 B3 B4 B5 B6 B7 gnd vdd
XNAND@0 A0 AB0 B0 gnd vdd NandGate_for8NAND__NAND
XNAND@1 A1 AB1 B1 gnd vdd NandGate_for8NAND__NAND
XNAND@2 A2 AB2 B2 gnd vdd NandGate_for8NAND__NAND
XNAND@3 A3 AB3 B3 gnd vdd NandGate_for8NAND__NAND
XNAND@4 A4 AB4 B4 gnd vdd NandGate_for8NAND__NAND
XNAND@5 A5 AB5 B5 gnd vdd NandGate_for8NAND__NAND
XNAND@6 A6 AB6 B6 gnd vdd NandGate_for8NAND__NAND
XNAND@7 A7 AB7 B7 gnd vdd NandGate_for8NAND__NAND
.ENDS _8Bit_NAND__8Bit_NAND

*** TOP LEVEL CELL: 8Bit_AND:8Bit_AND{lay}
X_8Bit_Inv@0 net@0 AandB0 net@2 AandB1 net@4 AandB2 net@6 AandB3 net@8 AandB4 net@10 AandB5 net@16 AandB6 net@14 AandB7 gnd vdd _8Bit_Inv__8Bit_Inv
X_8Bit_NAN@0 A0 A1 A2 A3 A4 A5 A6 A7 net@0 net@2 net@4 net@6 net@8 net@10 net@16 net@14 B0 B1 B2 B3 B4 B5 B6 B7 gnd vdd _8Bit_NAND__8Bit_NAND

* Spice Code nodes in cell cell '8Bit_AND:8Bit_AND{lay}'
vdd vdd 0 DC 5
va0 A0 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb0 B0 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va1 A1 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb1 B1 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va2 A2 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb2 B2 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va3 A3 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb3 B3 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va4 A4 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb4 B4 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va5 A5 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb5 B5 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va6 A6 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb6 B6 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va7 A7 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb7 B7 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.tran 200n
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
* Trailer cards described in this file:
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
.END
