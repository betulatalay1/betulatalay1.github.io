*** SPICE deck for cell left_shift{lay} from library left_shift
*** Created on Cum Ara 26, 2025 22:19:52
*** Last revised on Sal Ara 30, 2025 21:38:25
*** Written on Sal Ara 30, 2025 21:39:10 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Inverter_forleftshift__Inv FROM CELL Inverter_forleftshift:Inv{lay}
.SUBCKT Inverter_forleftshift__Inv gnd in out vdd
Mnmos@0 gnd in out gnd N L=0.6U W=3U AS=6.75P AD=18P PS=10.5U PD=28.5U
Mpmos@0 vdd in out vdd P L=0.6U W=3U AS=6.75P AD=20.25P PS=10.5U PD=29.1U
.ENDS Inverter_forleftshift__Inv

*** SUBCIRCUIT _8Bit_Inv_leftshift__8Bit_Inv FROM CELL 8Bit_Inv_leftshift:8Bit_Inv{lay}
.SUBCKT _8Bit_Inv_leftshift__8Bit_Inv A0 A1 A2 A3 A4 A5 A6 A7 gnd vdd Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
XInv@0 gnd A0 Y0 vdd Inverter_forleftshift__Inv
XInv@1 gnd A1 Y1 vdd Inverter_forleftshift__Inv
XInv@2 gnd A2 Y2 vdd Inverter_forleftshift__Inv
XInv@3 gnd A3 Y3 vdd Inverter_forleftshift__Inv
XInv@4 gnd A4 Y4 vdd Inverter_forleftshift__Inv
XInv@5 gnd A5 Y5 vdd Inverter_forleftshift__Inv
XInv@6 gnd A6 Y6 vdd Inverter_forleftshift__Inv
XInv@7 gnd A7 Y7 vdd Inverter_forleftshift__Inv
.ENDS _8Bit_Inv_leftshift__8Bit_Inv

*** SUBCIRCUIT buf_8__buf_8 FROM CELL buf_8:buf_8{lay}
.SUBCKT buf_8__buf_8 A0 A1 A2 A3 A4 A5 A6 A7 gnd vdd Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7
X_8Bit_Inv@0 A0 A1 A2 A3 A4 A5 A6 A7 gnd vdd net@45 net@34 net@30 net@27 net@23 net@20 net@17 net@14 _8Bit_Inv_leftshift__8Bit_Inv
X_8Bit_Inv@1 net@45 net@34 net@30 net@27 net@23 net@20 net@17 net@14 gnd vdd Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 _8Bit_Inv_leftshift__8Bit_Inv
.ENDS buf_8__buf_8

*** TOP LEVEL CELL: left_shift{lay}
Xbuf_8@0 gnd in0 in1 in2 in3 in4 in5 in6 gnd vdd Y0 Y1 Y2 Y3 Y4 Y5 Y6 Y7 buf_8__buf_8

* Spice Code nodes in cell cell 'left_shift{lay}'
vdd  vdd 0 DC 5
vin0 in0 0 DC pwl 10n 0 20n 5 50n 5 60n 0
vin1 in1 0 DC pwl 10n 0 20n 0 50n 0 60n 0
vin2 in2 0 DC pwl 10n 0 20n 5 50n 5 60n 0
vin3 in3 0 DC pwl 10n 0 20n 5 50n 5 60n 0
vin4 in4 0 DC pwl 10n 0 20n 0 50n 0 60n 0
vin5 in5 0 DC pwl 10n 0 20n 5 50n 5 60n 0
vin6 in6 0 DC pwl 10n 0 20n 0 50n 0 60n 0
vin7 in7 0 DC pwl 10n 0 20n 5 50n 5 60n 0
.tran 0 100ns
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
* Trailer cards described in this file:
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
.END
