*** SPICE deck for cell 8Bit_XOR{lay} from library 8Bit_XOR
*** Created on Sal Ara 23, 2025 21:42:40
*** Last revised on Sal Ara 23, 2025 22:08:38
*** Written on Sal Ara 23, 2025 22:08:41 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT XorGate_for8XOR__XOR FROM CELL XorGate_for8XOR:XOR{lay}
.SUBCKT XorGate_for8XOR__XOR A B gnd out vdd
Mnmos@0 net@6 A out gnd N L=0.6U W=3U AS=4.275P AD=5.4P PS=5.85U PD=8.1U
Mnmos@1 out net@17 net@6 gnd N L=0.6U W=3U AS=5.4P AD=4.275P PS=8.1U PD=5.85U
Mnmos@2 net@6 net@28 gnd gnd N L=0.6U W=3U AS=17.775P AD=5.4P PS=25.35U PD=8.1U
Mnmos@3 gnd B net@6 gnd N L=0.6U W=3U AS=5.4P AD=17.775P PS=8.1U PD=25.35U
Mnmos@4 gnd A net@28 gnd N L=0.6U W=3U AS=6.75P AD=17.775P PS=10.5U PD=25.35U
Mnmos@5 net@17 B gnd gnd N L=0.6U W=3U AS=17.775P AD=6.75P PS=25.35U PD=10.5U
Mpmos@0 vdd A net@1 vdd P L=0.6U W=3U AS=2.25P AD=21.6P PS=4.5U PD=27.9U
Mpmos@2 net@1 net@17 out vdd P L=0.6U W=3U AS=4.275P AD=2.25P PS=5.85U PD=4.5U
Mpmos@3 out net@28 net@4 vdd P L=0.6U W=3U AS=2.7P AD=4.275P PS=4.8U PD=5.85U
Mpmos@4 net@4 B vdd vdd P L=0.6U W=3U AS=21.6P AD=2.7P PS=27.9U PD=4.8U
Mpmos@5 vdd A net@28 vdd P L=0.6U W=3U AS=6.75P AD=21.6P PS=10.5U PD=27.9U
Mpmos@6 net@17 B vdd vdd P L=0.6U W=3U AS=21.6P AD=6.75P PS=27.9U PD=10.5U
.ENDS XorGate_for8XOR__XOR

*** TOP LEVEL CELL: 8Bit_XOR{lay}
XXOR@0 A0 B0 gnd AxorB_0 vdd XorGate_for8XOR__XOR
XXOR@1 A1 B1 gnd AxorB_1 vdd XorGate_for8XOR__XOR
XXOR@2 A2 B2 gnd AxorB_2 vdd XorGate_for8XOR__XOR
XXOR@3 A3 B3 gnd AxorB_3 vdd XorGate_for8XOR__XOR
XXOR@4 A4 B4 gnd AxorB_4 vdd XorGate_for8XOR__XOR
XXOR@5 A5 B5 gnd AxorB_5 vdd XorGate_for8XOR__XOR
XXOR@6 A6 B6 gnd AxorB_6 vdd XorGate_for8XOR__XOR
XXOR@7 A7 B7 gnd AxorB_7 vdd XorGate_for8XOR__XOR

* Spice Code nodes in cell cell '8Bit_XOR{lay}'
vdd vdd 0 DC 5
va0 A0 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb0 B0 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va1 A1 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb1 B1 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va2 A2 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb2 B2 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va3 A3 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb3 B3 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va4 A4 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb4 B4 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va5 A5 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb5 B5 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va6 A6 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb6 B6 0 DC pwl 10n 0 20n 5 100n 5 110n 0
va7 A7 0 DC pwl 10n 0 20n 5 50n 5 60n 0 90n 0 100n 5 130n 5 140n 0 170n 0 180n 5
vb7 B7 0 DC pwl 10n 0 20n 5 100n 5 110n 0
.tran 200n
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
* Trailer cards described in this file:
.include C:\Users\betul\OneDrive\Desktop\4-FALL\IC\C5_models.txt
.END
